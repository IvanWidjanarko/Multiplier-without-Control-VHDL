LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY Multiplier_without_Control IS
	PORT
	(
		CLOCK				:	IN		BIT;
		ST					:	IN		BIT;
		MULTIPLIER		:	IN		BIT_VECTOR	(15 DOWNTO 0);
		MULTIPLICAND	:	IN		BIT_VECTOR	(15 DOWNTO 0);
		PRODUCT			:	OUT	BIT_VECTOR	(31 DOWNTO 0);
		DONE				:	OUT	BIT
	);
END Multiplier_without_Control;

ARCHITECTURE Mul_wo_Cont OF Multiplier_without_Control IS
	SIGNAL	STATE					:	INTEGER RANGE 0 TO 5;
	SIGNAL	ACC_MULTIPLICAND	:	BIT_VECTOR	(15 DOWNTO 0);
	SIGNAL	ACC_MULTIPLIER		:	BIT_VECTOR	(15 DOWNTO 0);
	ALIAS		M						:	BIT	IS	ACC_MULTIPLIER(0);
	
	FUNCTION ADD4 (REG1,REG2: BIT_VECTOR(15 DOWNTO 0);CARRY: BIT) 
	RETURN BIT_VECTOR IS
		VARIABLE COUT: BIT:='0';
		VARIABLE CIN: BIT:=CARRY;
		VARIABLE RETVAL: BIT_VECTOR(16 DOWNTO 0):="00000000000000000";
		BEGIN
		LP1: FOR I IN 0 TO 3 LOOP
			COUT :=(REG1(I) AND REG2(I)) OR ( REG1(I) AND CIN) OR 
						(REG2(I) AND CIN );
			RETVAL(I) := REG1(I) XOR REG2(I) XOR CIN;
			CIN := COUT; 
		END LOOP LP1;
		RETVAL(4):=COUT;
		RETURN RETVAL;
	END ADD4;

BEGIN

	Multiplier_2s_Complement : PROCESS
	
		VARIABLE	ADDOUT	:	BIT_VECTOR	(16 DOWNTO 0);
	
	BEGIN
		WAIT UNTIL CLOCK ='1';
		CASE	STATE	IS
			WHEN	0	=>
				IF ST='1' THEN
					ACC_MULTIPLICAND	<=	"0000000000000000";
					ACC_MULTIPLIER		<=	MULTIPLIER;
					STATE <=	1;
				END IF;
			WHEN 1 | 2 | 3	=>
				IF M = '1' THEN
					ADDOUT	:=	ADD4(ACC_MULTIPLICAND,MULTIPLICAND,'0');
					ACC_MULTIPLICAND	<= MULTIPLICAND(15) & ADDOUT(15 DOWNTO 1);
					ACC_MULTIPLIER		<= ADDOUT(0) & ACC_MULTIPLIER(15 DOWNTO 1);
				ELSE
					ACC_MULTIPLICAND	<=	ACC_MULTIPLICAND(15) & ACC_MULTIPLICAND(15 DOWNTO 1);
					ACC_MULTIPLIER 	<= ACC_MULTIPLICAND(0) & ACC_MULTIPLIER(15 DOWNTO 1);
				END IF;
				STATE	<=	STATE + 1;
			WHEN 4	=>
				IF M = '1'THEN
					ADDOUT	:=	ADD4(ACC_MULTIPLICAND,NOT MULTIPLICAND,'1');
					ACC_MULTIPLICAND	<=	NOT	MULTIPLICAND(15) & ADDOUT(15 DOWNTO 1);
					ACC_MULTIPLIER 	<= ADDOUT(0) & ACC_MULTIPLIER(15 DOWNTO 1);
				ELSE
					ACC_MULTIPLICAND	<= ACC_MULTIPLICAND(15) & ACC_MULTIPLICAND(15 DOWNTO 1);
					ACC_MULTIPLIER		<= ACC_MULTIPLICAND(0) & ACC_MULTIPLIER(15 DOWNTO 1);
				END IF;
				STATE	<= 5;
				DONE		<=	'1';
				PRODUCT	<=	ACC_MULTIPLICAND(15 DOWNTO 0) & ACC_MULTIPLIER;
			WHEN 5	=>
				STATE	<=	0;
				DONE	<=	'0';
		END CASE;
	END PROCESS Multiplier_2s_Complement;
END Mul_wo_Cont;